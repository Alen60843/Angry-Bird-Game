//finish block background (remove white)

//finish random pig location

 

module houseMatrixBitMap(

	input logic clk,

	input logic resetN,

	input logic [10:0] offsetX,// offset from top left  position

	input logic [10:0] offsetY,

	input logic InsideRectangle, //input that the pixel is within a bracket

	input logic enterKey,

	input logic [4:0]randomX,

	input logic [4:0]randomY,

                                                                          
//------------------------input collision smiley and hart -student to complete functionality                                                                          

	input bird_house_collision,

	input bird_enemy_colision,

                                                                          

//------------------------random input

	input [21:0] randomHouse,

	input [8:0] randomPig_LVL,

	output  logic    drawingRequest, //output that the pixel should be dispalyed

	output logic fire,

	output  logic   [7:0] RGBout,  //rgb value from the bitmap
	
	output logic [10:0] pigLocationX,
	
	output logic [10:0] pigLocationY,

	output logic level1Vic,

	output logic level2Vic,

	output logic level3Vic,
	
	output logic preGame

) ;

 

 

// Size represented as Number of X and Y bits

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel

 /*  end generated by the tool */

 

 

// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 16*16 and use only the top left 16*15 squares

// this is the bitmap  of the maze , if there is a specific value  the  whole 32*32 rectange will be drawn on the screen

// there are  16 options of differents kinds of 32*32 squares

// all numbers here are hard coded to simplify the  understanding

 

enum logic [3:0] {PreGame,
	Idle,
	HouseLoad,
	PigDamageLoad,
	WinningScreen
	} SM_Motion;
 
logic enterKey_D;

logic level1;

logic level2;

logic level3;

logic currentLevel1;

logic currentLevel2;

logic currentLevel3;

logic currentLevel1_D;

logic currentLevel2_D;

logic currentLevel3_D;

logic enterKeyReg;

logic enterKeyReg_D;

logic enterKeyReg2;

logic enterKeyReg2_D;

logic bird_house_collision_D;

logic bird_enemy_colision_D;

 

int level;
int levelFlag;

 

logic [1:0] numOfPigs;

 

logic [0:15] [0:15] [3:0]  MazeBitMapMask ; 

 

logic [0:15] [0:15] [3:0]  defaultScreen= // level 1 option A

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000001234567800},

{64'h0000009ab0000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

logic [0:15] [0:15] [3:0]  MazeLVL1A= // level 1 option A

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000033300},

{64'h0000000000011100},

{64'h0000000000010100},

{64'h0000000003011100},

{64'h0000000001010101},// before 0000000001010100

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

 logic [0:15] [0:15] [3:0]  MazeLVL1B= // level 1 option B

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000030000000},

{64'h0000000010111110},

{64'h0000000010101010},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

 logic [0:15] [0:15] [3:0]  MazeLVL2A= // level 2 option A

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000083300},

{64'h0000000000015100},

{64'h0000000800050100},

{64'h0000000105151100},

{64'h0000000101010500},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

 logic [0:15] [0:15] [3:0]  MazeLVL2B= // level 2 option B

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000080000},

{64'h0000000301515100},

{64'h0000000101050100},

{64'h0000000505151100},

{64'h0000000101000500},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

 logic [0:15] [0:15] [3:0]  MazeLVL3A= // level 3 option A

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000888000},

{64'h0000000000555000},

{64'h0000000808505800},

{64'h0000000505555500},

{64'h0000000505050500},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

 logic [0:15] [0:15] [3:0]  MazeLVL3B= // level 3 option B

{{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000088800},

{64'h0000000003055500},

{64'h0000000801050500},

{64'h0000000505555500},

{64'h0000000505050500},

{64'h0000000000000000},

{64'h0000000000000000},

{64'h0000000000000000}};

 

//1 - wood square , 2 - wood square damaged, 3 - wood triangle , 4 - wood triangle damaged, 5 - stone square, 6 - stone square damaged mid , 7 - stone square damaged , 8 - stone triangle

//9 - stone triangle damaged mid , A - stone triangle damaged , B - pig

 

logic[0:10][0:31][0:31][7:0] object_colors = {
{	{8'hfa,8'hd5,8'hd1,8'hb1,8'hb1,8'hb0,8'hb0,8'hb0,8'hb0,8'hd0,8'hd0,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hb0,8'hb0,8'hb0,8'hb0,8'hb1,8'hd1,8'hd1,8'hd5,8'hda},
	{8'hb1,8'hd0,8'hf0,8'hf4,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hac},
	{8'hb0,8'hf5,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac},
	{8'hac,8'hf5,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hac,8'hf5,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'hac},
	{8'hac,8'hf5,8'hf4,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hac,8'hf5,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hcc,8'hf5,8'hf4,8'hf0,8'hf0,8'hf4,8'hf0,8'hd0,8'hd1,8'hd1,8'hd1,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd6,8'hfa,8'hfa,8'hda,8'hd5,8'hd5,8'hd5,8'hd5,8'hb1,8'hcc,8'hf0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac},
	{8'hcc,8'hf5,8'hf0,8'hf0,8'hf4,8'hf4,8'hd0,8'hfa,8'hfe,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf5,8'hf4,8'hf4,8'hf0,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf5,8'hf0,8'hf0,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hac,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf5,8'hf4,8'hf4,8'hf0,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf5,8'hf0,8'hf0,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf5,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hfe,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf5,8'hf0,8'hf0,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hcc,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hd0,8'hf5,8'hf0,8'hf0,8'hf0,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hd0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac},
	{8'hd0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hcc,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd5,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'h00,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfe,8'hfa,8'hd5,8'hac,8'hcc,8'hcc,8'hd0,8'hd0,8'hac,8'hac},
	{8'hcc,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hcc,8'hd0,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd1,8'hd5,8'hd1,8'hd1,8'hb1,8'hb1,8'hb1,8'hb1,8'hac,8'hac,8'hcc,8'hd0,8'hd0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac},
	{8'hac,8'hf9,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'hac},
	{8'hac,8'hf5,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hac,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hd0,8'hcc,8'hac,8'hac},
	{8'hac,8'hf5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac},
	{8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hcc,8'hac,8'hac,8'hac,8'hb1},
	{8'hd5,8'hac,8'hac,8'hac,8'hac,8'hcc,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'had,8'hd6}},

{	{8'hac,8'hac,8'hcc,8'hd0,8'hd0,8'hf1,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf5,8'hf5,8'hf5,8'hf0,8'hd0,8'hf0,8'hd0,8'hcc,8'hac,8'hac,8'h8c,8'h00},
	{8'hac,8'hf5,8'hf5,8'hf5,8'hf9,8'hf5,8'hf5,8'hf9,8'hf9,8'hf5,8'hf9,8'hf9,8'hf9,8'hf9,8'hf9,8'hf5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf5,8'hf9,8'hf9,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf5,8'hf0,8'hac,8'h00},
	{8'h00,8'h00,8'hd6,8'had,8'hac,8'hac,8'hac,8'hd0,8'hf1,8'hf5,8'hf5,8'hf5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf5,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hd1,8'hac,8'hac,8'hac,8'hac,8'hcc,8'hcc,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hd0,8'hd0,8'hd0,8'hf0,8'hd0,8'hac,8'hac,8'hfa},
	{8'hac,8'hd0,8'hf1,8'hf5,8'hf5,8'hf5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf5,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hfa},
	{8'hf5,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'hf6},
	{8'hf9,8'hf5,8'hf0,8'hf0,8'hf4,8'hf4,8'hf5,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hd5},
	{8'hf9,8'hf5,8'hf0,8'hf4,8'hf4,8'hf5,8'hac,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hd5},
	{8'hf5,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'had,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hac,8'hd1},
	{8'hf9,8'hf5,8'hf0,8'hf4,8'hf4,8'hf5,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hd1},
	{8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hd1},
	{8'hf9,8'hf4,8'hf0,8'hf0,8'hf4,8'hf1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'had,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hd6},
	{8'hf5,8'hf4,8'hf4,8'hf4,8'hf5,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf0,8'hf0,8'hd0,8'hac,8'hd5,8'h00,8'h00},
	{8'hf9,8'hf4,8'hf4,8'hac,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hac,8'hac,8'hac,8'hac,8'hac,8'h8c,8'hd1},
	{8'hf9,8'hf5,8'hd0,8'hf6,8'hac,8'hac,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'hd5},
	{8'hf5,8'hd0,8'hd0,8'hf4,8'hf4,8'hf1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'hd5},
	{8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'hd5},
	{8'hf9,8'hf5,8'hf4,8'hf4,8'hf4,8'hf1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hac,8'hac,8'hd1,8'hd0,8'hac,8'hac,8'hd6},
	{8'hf9,8'hf5,8'hf4,8'hf0,8'hf0,8'hd0,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'h00,8'hfa,8'hd1,8'hac,8'hac,8'hf6},
	{8'hd5,8'hf5,8'hac,8'hd0,8'hf0,8'hf1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb5,8'hac,8'hd0,8'hf0,8'hf0,8'hd0,8'hac,8'hfa},
	{8'hac,8'hd0,8'hf5,8'hf4,8'hf4,8'hf5,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'hfa},
	{8'hf9,8'hf9,8'hf4,8'hf4,8'hf4,8'hf5,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'hfe},
	{8'hf9,8'hf9,8'hf4,8'hf4,8'hf4,8'hf5,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'had,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hac,8'hfe},
	{8'hf9,8'hf9,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hcc,8'hcc,8'hcc,8'hcc,8'hac,8'hac,8'h00},
	{8'hf5,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hac,8'hac,8'hb1,8'hd6,8'hd6,8'hd6,8'hfa,8'hfa,8'h00,8'hfa,8'hfa,8'hd6,8'hd6,8'hd5,8'hb1,8'hac,8'hac,8'hac,8'hac,8'hd0,8'hd0,8'hf0,8'hf0,8'hcc,8'hac,8'h00},
	{8'hf9,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hac,8'h00},
	{8'hf5,8'hf9,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00},
	{8'hf5,8'hf5,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac,8'hd1,8'hb1,8'h8d,8'h00},
	{8'hf0,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'h00},
	{8'hcc,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hcc,8'hcc,8'hd0,8'hcc,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hf0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'hac,8'h00},
	{8'hac,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd5,8'h00},
	{8'had,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'had,8'hb1,8'hfa,8'h00,8'h00}},

 
 {	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hac,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf0,8'hf0,8'hac,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf0,8'hf0,8'hf0,8'hd0,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hf4,8'hf4,8'hf0,8'hcc,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hcc,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hcc,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hd0,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hd0,8'hf6,8'hd1,8'hf0,8'hf4,8'hf4,8'hf0,8'hf0,8'hac,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hd1,8'h00,8'hfa,8'hcc,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hcc,8'hfa,8'h00,8'h00,8'hd1,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hac,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hf0,8'hf4,8'hf0,8'hd1,8'h00,8'h00,8'h00,8'hfa,8'hd0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf0,8'hf4,8'hf4,8'hd0,8'hd0,8'hac,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hcc,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hac,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hfe,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hcc,8'hd0,8'hd0,8'hf0,8'hd0,8'hac,8'hd1,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd6,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'hd1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hfe,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf0,8'hf0,8'hf4,8'hf0,8'hd0,8'hd1,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'hd5,8'had,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hd1,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hd5,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf0,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hfa,8'h00,8'h00},
	{8'h00,8'h00,8'hd1,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hb1,8'h00,8'h00},
	{8'h00,8'hd5,8'hf5,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hfa,8'h00},
	{8'h00,8'hd1,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hf0,8'hd0,8'hac,8'hb1,8'h00},
	{8'hd5,8'hf5,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hfa},
	{8'hd0,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hd0,8'hd0,8'hf0,8'hf0,8'hf0,8'hd0,8'hcc,8'hac,8'hac,8'hac,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hb1},
	{8'hd0,8'hf5,8'hf0,8'hd0,8'hd0,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'hac,8'hac,8'hac,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'had},
	{8'hb1,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd6}},

 {	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfe,8'hac,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf4,8'hf4,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf4,8'hf0,8'hac,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hf5,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hcc,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hf0,8'hcc,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hac,8'hcc,8'hcc,8'hcc,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hd0,8'had,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'had,8'hac,8'hf5,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hcc,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf5,8'hf4,8'hf4,8'hf4,8'hf4,8'hcc,8'hf0,8'hd0,8'hf0,8'hf0,8'hf4,8'hd0,8'hd5,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hf9,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'hcc,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd0,8'hf5,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'h00,8'hac,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'hac,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf5,8'hac,8'h00,8'h00,8'hcc,8'hd0,8'hf0,8'hf0,8'hf4,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf5,8'hf4,8'hf4,8'hf0,8'hf0,8'hac,8'hfa,8'h00,8'h00,8'hac,8'hf5,8'hf4,8'hf4,8'hf4,8'hf5,8'hac,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hb1,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hfa,8'hd5,8'hd0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf0,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd1,8'hf5,8'hf4,8'hd0,8'hd0,8'hac,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd5,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hd0,8'hf0,8'hd0,8'hd0,8'hd0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hf9,8'hf4,8'hf4,8'hf4,8'hf4,8'hf5,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'had,8'hf5,8'hf0,8'hd0,8'hd0,8'hcc,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hfe,8'hf5,8'hf0,8'hf0,8'hf0,8'hf0,8'hf0,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hd0,8'hac,8'hac,8'hac,8'hac,8'h8c,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hac,8'hf4,8'hf4,8'hf4,8'hf4,8'hf4,8'hcc,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'had,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hb1,8'hf5,8'hd0,8'hf0,8'hf4,8'hf4,8'hf4,8'hac,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hac,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hac,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hf5,8'hf9,8'hf0,8'hf4,8'hf4,8'hf0,8'hf0,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hda,8'hf9,8'hf0,8'hf4,8'hf4,8'hf0,8'hf4,8'hf4,8'hf1,8'hd0,8'hf1,8'hf5,8'hf5,8'hf5,8'hf1,8'hd0,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hd0,8'hf4,8'hf4,8'hf0,8'hf4,8'hf4,8'hf0,8'hd0,8'hf0,8'hf4,8'hf4,8'hf0,8'hd0,8'hf0,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hac,8'h00,8'h00},
	{8'h00,8'h00,8'hf9,8'hf0,8'hf0,8'hf4,8'hf4,8'hd0,8'hac,8'hac,8'hf4,8'hf4,8'hf0,8'hf0,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hcc,8'hcc,8'hd0,8'hcc,8'hac,8'h00,8'h00},
	{8'h00,8'hac,8'hf5,8'hd0,8'hac,8'hac,8'hd1,8'hac,8'hf5,8'hf4,8'hd0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'had,8'h00},
	{8'h8d,8'h8c,8'hb1,8'h00,8'h00,8'hf6,8'hac,8'hf5,8'hd0,8'hf0,8'hf4,8'hf4,8'hf4,8'hf0,8'hd0,8'hd0,8'hcc,8'hd0,8'hcc,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hcc,8'hac,8'hd6},
	{8'h00,8'h00,8'h00,8'h00,8'hfa,8'hac,8'hd0,8'hcc,8'hd0,8'hf0,8'hf0,8'hf0,8'hd0,8'hac,8'hac,8'hf5,8'hac,8'hcc,8'hcc,8'hd0,8'hcc,8'hcc,8'hcc,8'hd0,8'hcc,8'hd0,8'hd0,8'hac,8'hac,8'hac,8'hac,8'h8c},
	{8'h00,8'h00,8'h00,8'hac,8'hcc,8'hac,8'hd0,8'hd0,8'hd0,8'hd0,8'hd0,8'hac,8'hfa,8'hf5,8'hf5,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hcc,8'hac,8'hac,8'hac,8'hac,8'hac,8'hcc,8'hcc,8'hac,8'h8c},
	{8'h00,8'h00,8'h8d,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hd6,8'h8c,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hac,8'hb1}},

 
{	{8'hb6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h92},
	{8'h6d,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hfb,8'hb2,8'h6d},
	{8'h6d,8'h00,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'hd6,8'hd6,8'hd6,8'hb2,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'h00,8'hd6,8'hb6,8'hb1,8'hb1,8'hb1,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'hfb,8'hb1,8'hb1,8'hb6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb6,8'hb6,8'hb2,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h8d,8'h8d,8'h91,8'h91,8'h91,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'h91,8'h00,8'hb6,8'hd6,8'hd6,8'hd6,8'h8d,8'h91,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hb2,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'hb2,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hb6,8'hb1,8'h8d,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb6,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb2,8'hb1,8'hb1,8'h91,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hd6,8'hfb,8'hb2,8'h8d,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb6,8'hb2,8'hb1,8'h91,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb2,8'hb1,8'hb1,8'h91,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb1,8'hb1,8'hb1,8'h91,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'hb2,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h6d,8'h8d,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb2,8'h91,8'h91,8'h8d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h8d,8'h6d,8'h8d,8'h91,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'h00,8'hd6,8'hd6,8'h91,8'h91,8'hd6,8'hb6,8'hb1,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'hfb,8'hb2,8'hb1,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h8d,8'h6d},
	{8'h6d,8'hfb,8'hb1,8'hb1,8'hb2,8'hfb,8'hd6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h8d,8'h6d},
	{8'h6d,8'hfb,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h8d,8'h6d,8'h6d},
	{8'h6d,8'h6d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h91,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h6d,8'h6d,8'h6d,8'h6d,8'h92},
	{8'hd6,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'hb6,8'h00,8'h00}},
 
  
 {	{8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h65,8'h00},
	{8'h24,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfb,8'hb6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h6d,8'h6d},
	{8'h91,8'hff,8'hda,8'hb6,8'hb6,8'hb6,8'hb6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'h91,8'h8d,8'h91,8'hd6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb1,8'h6d,8'h6d,8'h24},
	{8'hb6,8'hff,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'h8d,8'h8d,8'h91,8'hd6,8'hb6,8'hd6,8'h8d,8'hb6,8'hd6,8'hd6,8'hd6,8'hb1,8'h8d,8'h8d,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h00,8'hd6,8'h8d,8'hb6,8'hd6,8'hb1,8'h91,8'h91,8'h24},
	{8'hff,8'hff,8'hd6,8'hb1,8'h91,8'h91,8'hb1,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h91,8'h91,8'h24},
	{8'hff,8'hd6,8'hb1,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'hda,8'hb6,8'hb1,8'h91,8'h91,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'h8d,8'hb1,8'h91,8'h91,8'h24},
	{8'hff,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'h24,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hd6,8'hd6,8'hb6,8'hd6,8'h91,8'h91,8'h24},
	{8'hff,8'hda,8'hd6,8'hd6,8'hd6,8'hda,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'hd6,8'hd6,8'hd6,8'h91,8'h91,8'h91,8'h25},
	{8'hb1,8'h91,8'hd6,8'hd6,8'hd6,8'hb6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hda,8'hd6,8'hd6,8'h8d,8'hb1,8'h91,8'h25},
	{8'hff,8'h8d,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'hd6,8'h8d,8'hb2,8'h91,8'h25},
	{8'hff,8'hda,8'h8d,8'h91,8'h8d,8'h91,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'hd6,8'h8d,8'hb2,8'h91,8'h25},
	{8'hff,8'hda,8'hd6,8'h8d,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'hd6,8'h8d,8'hb6,8'h91,8'h25},
	{8'hff,8'hda,8'hd6,8'hb1,8'hd6,8'hb6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb2,8'hd6,8'hd6,8'h8d,8'hb6,8'h91,8'h25},
	{8'hff,8'hda,8'hd6,8'hd6,8'hd6,8'hb2,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'hb6,8'h91,8'hb6,8'h91,8'h65},
	{8'hff,8'hda,8'hb6,8'hd6,8'hb6,8'hb6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'hd6,8'hda,8'h91,8'hb6,8'h91,8'h24},
	{8'hff,8'hda,8'hd6,8'hd6,8'h91,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h8d,8'h00,8'hfb,8'hb6,8'h91,8'h24},
	{8'hff,8'hda,8'hd6,8'hd6,8'h8d,8'hb6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'h91,8'hb2,8'hb6,8'h91,8'h24},
	{8'hff,8'hfa,8'hd6,8'hd6,8'hb1,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'hb1,8'hb2,8'hb6,8'h91,8'h24},
	{8'hff,8'hfb,8'hd6,8'hd6,8'hb6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb6,8'hb2,8'hb2,8'hb2,8'h91,8'h24},
	{8'hff,8'hfb,8'hd6,8'hd6,8'hd6,8'hd6,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb1,8'hb2,8'h91,8'hb6,8'h91,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'h91,8'hd6,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb1,8'hb1,8'h91,8'hb6,8'h91,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'hd6,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb2,8'hb1,8'h8d,8'hb1,8'h91,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'h8d,8'hda,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hb6,8'hb1,8'hb1,8'h91,8'h91,8'h8d,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'hb1,8'hda,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h24,8'hb6,8'hb1,8'hb2,8'h91,8'hb1,8'h8d,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'hd6,8'hb2,8'hda,8'hb6,8'hb2,8'h91,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h6d,8'h6d,8'h8d,8'hb1,8'hb6,8'hb6,8'hb2,8'hb1,8'hb1,8'hb1,8'h91,8'hb1,8'h6d,8'h24},
	{8'hff,8'hff,8'hd6,8'hd6,8'h8d,8'h8d,8'hb6,8'h8d,8'h91,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'hb2,8'h91,8'h6d,8'h6d},
	{8'hfb,8'hff,8'hb2,8'h8d,8'hd6,8'hd6,8'hd6,8'h8d,8'hd6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb2,8'hb1,8'hb2,8'h91,8'h91,8'h8d,8'h8d,8'h91,8'h91,8'h91,8'hb1,8'h8d,8'h6d,8'h91},
	{8'hb6,8'hff,8'h91,8'h91,8'hd6,8'h00,8'h91,8'hb2,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb2,8'h91,8'hb1,8'hb2,8'hb2,8'h8d,8'h91,8'h91,8'hb1,8'hb1,8'hb2,8'h8d,8'h6d,8'hda},
	{8'h6d,8'hff,8'h91,8'hb1,8'hb2,8'hb6,8'hb2,8'hb2,8'hb2,8'h91,8'hb2,8'hb2,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb2,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb2,8'h91,8'hb2,8'hb6,8'h91,8'h8d,8'h8d,8'h6d,8'h00},
	{8'h65,8'h6d,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h8d,8'h91,8'h91,8'h8d,8'h8d,8'h8d,8'h8d,8'h8d,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h8d,8'h6d,8'h6d,8'h6d,8'h24,8'h00},
	{8'h24,8'h24,8'h25,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24,8'h24,8'h24,8'h6d,8'hb6,8'h00,8'h00}},

	
{	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h24},
	{8'h00,8'h00,8'h00,8'h91,8'h91,8'hb6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'h20,8'h00,8'h00,8'hda,8'h8d,8'h64,8'h6d,8'h00,8'hd6,8'hb6,8'hb6,8'hd6,8'h91,8'hb6,8'h91,8'h24},
	{8'h00,8'h00,8'hb2,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h24,8'h00,8'h00,8'h91,8'hd6,8'h6d,8'h24,8'h00,8'hb2,8'hd6,8'hb1,8'hd6,8'h91,8'h24},
	{8'h00,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'h64,8'h91,8'h00,8'hfb,8'hb6,8'hb1,8'hb2,8'hb6,8'h91,8'h91,8'h00,8'h64,8'h24,8'h00,8'h91,8'hb6,8'h8d,8'h24},
	{8'h00,8'h00,8'hda,8'hb6,8'h8d,8'h6d,8'h6d,8'hb6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hd6,8'hd6,8'hb6,8'hb6,8'hb6,8'hd6,8'hb1,8'h8d,8'hb6,8'hd6,8'h00,8'h00,8'hb6,8'hb6,8'h6d,8'h65},
	{8'h00,8'h00,8'h91,8'h91,8'hda,8'hd6,8'hd6,8'hfa,8'h00,8'h00,8'hfb,8'hda,8'hb6,8'h8d,8'h91,8'h91,8'h65,8'h65,8'h6c,8'h64,8'h6d,8'h91,8'h6d,8'hb6,8'hda,8'hda,8'hd6,8'h65,8'h00,8'hb6,8'h00,8'h00},
	{8'h00,8'h00,8'hda,8'hb6,8'hd6,8'hb6,8'h24,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hb6,8'hfb,8'h64,8'h24,8'h00,8'h24},
	{8'h00,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb6,8'hd6,8'h6d,8'h24,8'h24,8'h65},
	{8'hb6,8'h00,8'h00,8'hb6,8'hd6,8'hd6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb6,8'h24,8'hda,8'h91,8'h6d},
	{8'h91,8'h00,8'h24,8'h00,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'h64,8'h91,8'h91,8'h6d},
	{8'hb2,8'h00,8'h6d,8'h6d,8'h24,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hd6,8'hb6,8'h00,8'h91,8'h6d},
	{8'hb6,8'h00,8'hd6,8'hda,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'h8d,8'h00,8'h91,8'h6d},
	{8'hb6,8'h00,8'hd6,8'h00,8'h24,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'h24,8'h6d,8'h91,8'h6d},
	{8'hd6,8'h00,8'hd6,8'hda,8'h6d,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'h6d,8'h00,8'h91,8'h6d},
	{8'hda,8'h00,8'hd6,8'hd6,8'h6d,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h6d,8'h00,8'h91,8'h6d},
	{8'hda,8'h00,8'hd6,8'hd6,8'h24,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'h6d,8'h00,8'hda,8'h91,8'h65},
	{8'hda,8'h00,8'hd6,8'hd6,8'h24,8'hfa,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h24,8'h00,8'h6d,8'h8d,8'h65},
	{8'hda,8'h00,8'hd6,8'hb6,8'h24,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hb1,8'h00,8'h8d,8'h8d,8'h24},
	{8'hb6,8'h00,8'hd6,8'hd6,8'h24,8'hb6,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb2,8'h00,8'hd6,8'h8d,8'h24},
	{8'hb6,8'h00,8'hd6,8'hda,8'h24,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb1,8'h24,8'h00,8'h8d,8'h24},
	{8'hb5,8'h00,8'hd6,8'hfb,8'h91,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb1,8'h6d,8'h00,8'h6d,8'h24},
	{8'h91,8'h00,8'hd6,8'hda,8'h20,8'h24,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb6,8'hb1,8'h6d,8'h00,8'h24,8'h00},
	{8'h6d,8'h00,8'hd6,8'hb6,8'h24,8'h00,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hb1,8'hb1,8'h64,8'h6d,8'h00,8'h24},
	{8'h24,8'h00,8'hd6,8'hd6,8'hb1,8'hfb,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h00,8'h24,8'hb1,8'hb2,8'h6d,8'h00,8'h64,8'h25},
	{8'h00,8'h00,8'hd6,8'hd6,8'hfa,8'h24,8'h00,8'h00,8'hd6,8'h8d,8'h6d,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6c,8'h6c,8'h6d,8'h91,8'hd6,8'hda,8'hb6,8'hb1,8'hb2,8'hb6,8'h24,8'h00,8'h91,8'h24},
	{8'h00,8'h00,8'hd6,8'hd6,8'h6d,8'h8d,8'h24,8'h00,8'h24,8'hd6,8'hd6,8'hb6,8'hb6,8'hd6,8'hb6,8'hb6,8'hd6,8'hda,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb2,8'hb6,8'h6d,8'hda,8'h91,8'h91,8'h24},
	{8'h00,8'h00,8'hb1,8'h24,8'h04,8'h00,8'h00,8'h24,8'hb1,8'h00,8'hd6,8'hd6,8'hd6,8'hda,8'hb2,8'h91,8'hb1,8'hb1,8'hb2,8'hb1,8'hb6,8'hb1,8'h6d,8'h64,8'h64,8'h00,8'hb6,8'h24,8'h91,8'hd6,8'h91,8'h00},
	{8'h00,8'h00,8'hb2,8'h6d,8'hb2,8'h00,8'hda,8'hb1,8'hd6,8'h24,8'h00,8'hb2,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb6,8'hb6,8'h24,8'hda,8'h00,8'h24,8'h00,8'h8d,8'h00,8'hfa,8'hb2,8'h91,8'h91,8'h00},
	{8'h04,8'h00,8'h91,8'h24,8'hb2,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb6,8'h24,8'h6d,8'hd6,8'hb1,8'hb1,8'hb2,8'h91,8'h65,8'h00,8'hb1,8'h6d,8'h8d,8'h6d,8'h00},
	{8'h00,8'h20,8'h91,8'h24,8'h24,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'h00,8'h8d,8'h8d,8'h8d,8'h8d,8'h65,8'h24,8'hda,8'h65,8'h8d,8'h91,8'h91,8'h8d,8'h00,8'hb2,8'h91,8'h6d,8'h6d,8'h64,8'h6d,8'h00},
	{8'hb2,8'h00,8'h00,8'h24,8'h24,8'h24,8'h65,8'h24,8'h24,8'h64,8'h64,8'h00,8'h24,8'h24,8'h24,8'h24,8'h24,8'h00,8'h24,8'h24,8'h25,8'h24,8'h25,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'h00}},

	
{	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hd6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h00,8'hd6,8'hd6,8'hb2,8'hb2,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hda,8'hd6,8'hd6,8'hd6,8'hb6,8'h8d,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'hb2,8'hd6,8'hd6,8'hb2,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hb1,8'hd6,8'hb1,8'hd6,8'hd6,8'hb2,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'hd6,8'hd6,8'hd6,8'hb1,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hb2,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hfb,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h00,8'hda,8'hb1,8'hd6,8'hd6,8'hb6,8'h6d,8'h91,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hb6,8'hd6,8'hd6,8'hb2,8'h91,8'h6d,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hfb,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h8d,8'hb2,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h91,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb2,8'h91,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb2,8'hd6,8'hd6,8'hd6,8'hd6,8'hb2,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'hd6,8'hd6,8'hb6,8'h91,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'hd6,8'hb2,8'hb1,8'h91,8'hb6,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h91,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'hda,8'hb1,8'hb1,8'h91,8'h6d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hb2,8'hb1,8'hb1,8'hb1,8'h8d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb2,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hb6,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hb6,8'hda,8'hda,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h6d,8'h91,8'h00,8'h00},
	{8'h00,8'h00,8'hb6,8'h00,8'hd6,8'hd6,8'h91,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'hb2,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hda,8'hb2,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h8d,8'hb6,8'h00},
	{8'h00,8'h8d,8'h00,8'hd6,8'hd6,8'hd6,8'hda,8'hfa,8'hfa,8'hd6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h6d,8'h00},
	{8'h6d,8'hfb,8'hb2,8'hb1,8'hb1,8'hb6,8'hb6,8'hb6,8'hb6,8'hd6,8'hda,8'hda,8'hb6,8'hb6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h91,8'h6d},
	{8'h8d,8'h00,8'hb1,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h8d,8'hfb,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d}},

	
{	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h6d,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hda,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hb6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h00,8'hd6,8'h91,8'hb1,8'hb2,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hb6,8'hb2,8'hd6,8'hb6,8'hb6,8'h8d,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'hb6,8'h91,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hb6,8'h91,8'hd6,8'hd6,8'hb2,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hb1,8'h91,8'hb1,8'hd6,8'hd6,8'hb2,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'hd6,8'hd6,8'hd6,8'h91,8'hd6,8'hd6,8'hd6,8'hb6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hd6,8'hb1,8'hb6,8'hda,8'hd6,8'hd6,8'hd6,8'hb1,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'hb2,8'hda,8'hd6,8'hb6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hfb,8'hd6,8'hb1,8'hb6,8'hd6,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfb,8'h00,8'hda,8'h91,8'hb6,8'hd6,8'hb6,8'h6d,8'h91,8'hd6,8'hd6,8'hd6,8'hb1,8'hb6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'h91,8'hd6,8'hd6,8'hb2,8'h91,8'h6d,8'hb6,8'hd6,8'hd6,8'h91,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hfb,8'hd6,8'hb6,8'hb6,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'h91,8'hd6,8'hd6,8'h8d,8'hb2,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'h00,8'hd6,8'hb6,8'hd6,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h91,8'hb6,8'hd6,8'h91,8'hd6,8'hd6,8'hb1,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hda,8'h00,8'hd6,8'hd6,8'h91,8'hd6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h91,8'hb1,8'hb6,8'hd6,8'hb6,8'h91,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hb6,8'h91,8'hd6,8'hb2,8'h91,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb2,8'hd6,8'h91,8'hd6,8'hd6,8'hb2,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'h91,8'hb2,8'hb6,8'hb6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'h91,8'hd6,8'hd6,8'h6d,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h00,8'hd6,8'hd6,8'h91,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'hb6,8'hb2,8'hb6,8'h91,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hd6,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hd6,8'hd6,8'h91,8'h91,8'hb1,8'h91,8'hb6,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h91,8'hda,8'hd6,8'hd6,8'hb6,8'hd6,8'hb6,8'hda,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'h91,8'hda,8'hb1,8'hb1,8'h91,8'h6d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'hd6,8'hd6,8'hd6,8'hb6,8'hd6,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hb6,8'hb2,8'hb1,8'h91,8'hb1,8'h8d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h6d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'hb1,8'hb1,8'hb1,8'h91,8'h91,8'h6d,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'hb6,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hb6,8'hb6,8'hb6,8'hb6,8'h91,8'h91,8'hb6,8'hb6,8'hda,8'hda,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'hb1,8'h6d,8'h91,8'h00,8'h00},
	{8'h00,8'h00,8'hb6,8'h00,8'hd6,8'hd6,8'h91,8'h91,8'hb6,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hb6,8'hd6,8'hda,8'hb2,8'hb1,8'h91,8'hb1,8'hb1,8'hb1,8'h91,8'h91,8'hb1,8'h91,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hb1,8'hb1,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'h91,8'hb6,8'hb2,8'hb1,8'hb1,8'h91,8'hb1,8'hb1,8'hb1,8'h91,8'hb1,8'hb1,8'h91,8'h8d,8'hb6,8'h00},
	{8'h00,8'h8d,8'h00,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h91,8'hb2,8'h91,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb1,8'hb1,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'hb1,8'hb1,8'hb1,8'h91,8'h6d,8'h00},
	{8'h6d,8'hfb,8'hb2,8'hb1,8'hb1,8'h91,8'hb1,8'hb6,8'hd6,8'hd6,8'hda,8'hda,8'hb6,8'hb6,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'hb1,8'h91,8'h91,8'h6d},
	{8'h8d,8'h00,8'hb1,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h8d,8'hfb,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d}},

	
{	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hfa,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hb6,8'h6d,8'hb6,8'h91,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hb6,8'h6d,8'hda,8'h91,8'hd6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'hff,8'h6d,8'hda,8'hd6,8'hb2,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hda,8'hd6,8'h6d,8'hd6,8'hd6,8'hb1,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hff,8'hb6,8'h91,8'h6d,8'hb1,8'hd6,8'hd6,8'hb1,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hb6,8'hd6,8'hd6,8'h8d,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'hff,8'hd6,8'hd6,8'h91,8'h6d,8'hfa,8'hb6,8'hd6,8'hd6,8'hb6,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h91,8'hd6,8'hd6,8'hd6,8'h6d,8'hfb,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h65,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hd6,8'h91,8'h6d,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hda,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hd6,8'h8d,8'hb6,8'hd6,8'hd6,8'h24,8'h91,8'hd6,8'hd6,8'hb6,8'h91,8'hda,8'hb1,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hb6,8'h6d,8'hd6,8'hb6,8'hb6,8'h6d,8'h24,8'hda,8'hd6,8'hd6,8'h91,8'hd6,8'hb1,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'hb6,8'hd6,8'h8d,8'hd6,8'hd6,8'h24,8'h00,8'h00,8'h24,8'hd6,8'hd6,8'h6d,8'hb6,8'hd6,8'h6d,8'h8d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hff,8'hd6,8'hb6,8'hfb,8'hd6,8'hda,8'hfb,8'h00,8'h00,8'h8d,8'hd6,8'hd6,8'h6d,8'hb6,8'hd6,8'hb2,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hdb,8'hff,8'hb6,8'hd6,8'h6d,8'hda,8'hd6,8'h24,8'h00,8'h00,8'h00,8'h00,8'h24,8'h6d,8'h6d,8'hd6,8'hb6,8'hd6,8'hb1,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hff,8'hd6,8'hda,8'h6d,8'hb6,8'hb6,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h65,8'hb6,8'hd6,8'h6d,8'hfb,8'hd6,8'hb2,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h65,8'h6d,8'h6d,8'hb6,8'h91,8'hb2,8'hd6,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hd6,8'hd6,8'h6d,8'hd6,8'hd6,8'h6d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hff,8'hb6,8'hb6,8'h6d,8'h00,8'hd6,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb6,8'hd6,8'h91,8'hb2,8'hb6,8'h91,8'h64,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hb6,8'hff,8'hb6,8'hd6,8'hd6,8'h6d,8'hd6,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'hd6,8'hd6,8'h6d,8'h91,8'hb1,8'h91,8'hb2,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h6d,8'hda,8'hd6,8'hd6,8'h8d,8'h00,8'hd6,8'hfb,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'hb1,8'h6d,8'h00,8'h8d,8'h00,8'h91,8'h65,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hff,8'hb6,8'hd6,8'hd6,8'h6d,8'h00,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h91,8'hb1,8'hb2,8'h6d,8'hfb,8'h6d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'hff,8'hd6,8'hd6,8'hd6,8'hb6,8'h91,8'h24,8'h20,8'h00,8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h24,8'h65,8'hb1,8'hb1,8'h91,8'h6d,8'h91,8'h24,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h91,8'hff,8'hb6,8'hd6,8'hd6,8'hd6,8'hd6,8'h6d,8'h00,8'hda,8'hda,8'hda,8'h8d,8'h91,8'h00,8'h00,8'h00,8'h00,8'h6d,8'h00,8'hb6,8'hb2,8'hb1,8'hb2,8'h6d,8'hb6,8'h6d,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'hb2,8'hff,8'hb6,8'hd6,8'h91,8'h91,8'hd6,8'h6d,8'hfa,8'hd6,8'hd6,8'hd6,8'hd6,8'h8d,8'hfb,8'hd6,8'hfb,8'hb1,8'hb2,8'h6d,8'hfa,8'hb1,8'hb1,8'h6d,8'hb6,8'hb1,8'h91,8'h6d,8'h00,8'h00},
	{8'h00,8'h00,8'hff,8'hda,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'h6d,8'h8d,8'hb6,8'hd6,8'hd6,8'hb6,8'hd6,8'h6d,8'h91,8'h91,8'hb6,8'hb6,8'h6d,8'hd6,8'hb6,8'hb6,8'h6d,8'h00,8'hb1,8'h91,8'h8d,8'hb6,8'h00},
	{8'h00,8'h24,8'hff,8'hd6,8'hd6,8'hd6,8'hda,8'h6d,8'h6d,8'hb6,8'h6d,8'hd6,8'hd6,8'hd6,8'hd6,8'hb6,8'hfa,8'hb1,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h91,8'h91,8'hb1,8'hb2,8'h91,8'h65,8'h00},
	{8'h24,8'hff,8'h91,8'hb2,8'hb2,8'h65,8'hb6,8'hfa,8'hd6,8'hd6,8'h00,8'h00,8'hb6,8'hb2,8'hb1,8'hb1,8'hb1,8'hb1,8'hb6,8'h6d,8'hd6,8'h91,8'h91,8'h91,8'h91,8'hb1,8'hb2,8'hb2,8'hb2,8'h91,8'h91,8'h24},
	{8'h24,8'hff,8'hb2,8'h91,8'h6d,8'hd6,8'h8d,8'h8d,8'h8d,8'h91,8'h8d,8'h6d,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h6d,8'h00,8'h91,8'h91,8'h91,8'h91,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h6d,8'hff,8'h91,8'h8d,8'h00,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h8d,8'hb6,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d,8'hfb,8'h8d,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h91,8'h6d},
	{8'h24,8'h24,8'h6d,8'h6d,8'h24,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h64,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h65,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h6d,8'h24}},

	
{	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h9d,8'h9d,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h04,8'h04,8'h9d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h99,8'h9d,8'h9d,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h04,8'h04,8'h9d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h74,8'h04,8'h9d,8'h00,8'h00,8'h00,8'h2c,8'h30,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h30,8'h04,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'hbd,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'hbd,8'hbd,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'hbd,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'h74,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h2c,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'hbd,8'h0c,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h9d,8'h9d,8'h78,8'h9c,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h34,8'h9d,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h9d,8'h9d,8'h30,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h7c,8'h78,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h78,8'h74,8'h74,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h74,8'h00,8'h00},
	{8'h00,8'h04,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h98,8'hdc,8'hdc,8'hdc,8'hdc,8'hbc,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h00,8'h00},
	{8'h00,8'h7c,8'h9d,8'h9d,8'h9d,8'h74,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'hbc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hfc,8'hfc,8'hdc,8'h9c,8'h9d,8'h9d,8'h9d,8'h74,8'h95,8'h95,8'h9c,8'h9d,8'h00,8'h00},
	{8'h00,8'h9d,8'h9d,8'h9d,8'h95,8'hff,8'hff,8'hba,8'h9d,8'h9d,8'h74,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hfc,8'hbc,8'h9d,8'h9d,8'h78,8'hff,8'hff,8'hff,8'hff,8'h78,8'h30,8'h00},
	{8'h00,8'h9d,8'h78,8'hb9,8'hff,8'hff,8'hff,8'hff,8'hff,8'h74,8'hdc,8'hdc,8'hdc,8'h04,8'h04,8'hdc,8'hdc,8'hdc,8'hb8,8'hdc,8'hdc,8'hdc,8'h98,8'h78,8'hde,8'hff,8'hff,8'hda,8'hff,8'hff,8'h9d,8'h00},
	{8'h00,8'h9d,8'h78,8'hff,8'hff,8'h00,8'hb6,8'hff,8'hff,8'h98,8'hdc,8'hdc,8'h70,8'h04,8'h04,8'h70,8'hdc,8'hdc,8'h04,8'h04,8'hdc,8'hfc,8'hdc,8'h78,8'hff,8'hff,8'hff,8'hda,8'hff,8'hff,8'h9d,8'h00},
	{8'h00,8'h9d,8'h78,8'hde,8'hff,8'hb6,8'hff,8'hff,8'hff,8'hbc,8'hdc,8'hdc,8'h30,8'h04,8'h04,8'h2c,8'hdc,8'hbc,8'h04,8'h04,8'hdc,8'hdc,8'hdc,8'h78,8'hda,8'hff,8'hff,8'hff,8'hff,8'hff,8'h9d,8'h00},
	{8'h00,8'h9c,8'h78,8'h70,8'hff,8'hff,8'hff,8'hff,8'h74,8'h98,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'h78,8'h74,8'hff,8'hff,8'hff,8'hda,8'h78,8'h9c,8'h00},
	{8'h00,8'h7c,8'h9d,8'h78,8'h70,8'h95,8'hb5,8'h70,8'h9d,8'h74,8'hbc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'h9d,8'h78,8'h70,8'h70,8'h70,8'h78,8'h9d,8'h7c,8'h00},
	{8'h00,8'h30,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h98,8'hbc,8'hbc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hdc,8'hbc,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h04,8'h00},
	{8'h00,8'h00,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h74,8'h98,8'h98,8'hb8,8'hbc,8'hbc,8'hbc,8'hbc,8'h98,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h00,8'h00},
	{8'h00,8'h00,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h74,8'h98,8'h98,8'h98,8'h98,8'h98,8'h98,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h78,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h94,8'h98,8'h98,8'h98,8'h74,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h78,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h78,8'h78,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h78,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h78,8'h7c,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h7c,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h78,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h78,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h78,8'h7c,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9d,8'h9c,8'h78,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h34,8'h78,8'h78,8'h78,8'h78,8'h78,8'h34,8'h30,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
	{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}
	}};


// assign offsetY_LSB  = offsetY[4:0] ; // get lower 5 bits

// assign offsetY_MSB  = offsetY[8:5] ; // get higher 4 bits

// assign offsetX_LSB  = offsetX[4:0] ;

// assign offsetX_MSB  = offsetX[8:5] ;

 

// pipeline (ff) to get the pixel color from the array           

 

//==----------------------------------------------------------------------------------------------------------------=

always_ff@(posedge clk or negedge resetN)

begin

	if(!resetN) begin

		RGBout <=         8'h00;

		MazeBitMapMask  <=  defaultScreen;  //  copy default tabel

		enterKey_D <= 0; //remembers enter after 1 cycle

		level1Vic <= 0;

		level2Vic <= 0;

		level3Vic <= 0;

		levelFlag <= 0;
		
		preGame <= 1;

		level <= 1;
		
		SM_Motion <= PreGame;


	end

	else begin
	
		case(SM_Motion)
		
			//--------

				PreGame: begin

			//--------
				enterKey_D <= enterKey;
				if(enterKey && !enterKey_D) begin
					SM_Motion <= Idle;
					preGame <= 0;
				end
			
			end

			//--------

				Idle: begin

			//--------

					enterKey_D <= enterKey;

					if(levelFlag == 0)

						SM_Motion <= HouseLoad;

																	  

                                            

					RGBout <= TRANSPARENT_ENCODING ; // default

					bird_house_collision_D <= bird_house_collision;

					bird_enemy_colision_D <= bird_enemy_colision;

                                            

////////////////////////////////////////////////////////colision

					if (bird_house_collision && !bird_house_collision_D)begin

						if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h1 ) //wood square to damaged wood square

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h2;

						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h2)     //damaged wood squared destroyed

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;

						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h3) // wood triangle to damaged wood triangle

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h4;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h4) // wood triangle damaged destroyed

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h5) // stone square to stone square damaged mid

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h6;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h6) // stone square damaged mid to stone square damaged

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h7;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h7) // stone square damaged destroyed

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;
								

						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h8) // stone triangle to stone triangle damaged mid

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h9;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'h9) // stone triangle damaged mid to stone triangle damaged

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'hA;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'ha) // stone triangle damaged destroyed

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;


						else if(MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] == 4'hb) begin // pig destroyed

								MazeBitMapMask[offsetY[8:5]][offsetX[8:5]] <= 4'h0;

								if(level == 1) begin

									level <= 2;

									level1Vic <= 1;
									
									SM_Motion <= WinningScreen;

									end

								else if (level == 2) begin

									level <= 3;

									level2Vic <= 1;
									
									SM_Motion <= WinningScreen;

									end

								else if (level == 3) begin

									level <= 1;

									level3Vic <= 1;
									
									SM_Motion <= WinningScreen;

									end


								end

                                                           

						end

                                                                          

                                                                                                        

////////////////////////////////////////////////////////

					if (InsideRectangle == 1'b1 )     

						begin

							case (MazeBitMapMask[offsetY[8:5]][offsetX[8:5]])

								4'h0 : RGBout <= TRANSPARENT_ENCODING ;

								4'h1 : RGBout <= object_colors[4'h0][offsetY[4:0]][offsetX[4:0]]; // wood square

								4'h2 : RGBout <= object_colors[4'h1][offsetY[4:0]][offsetX[4:0]] ;// wood square damaged

								4'h3 : RGBout <= object_colors[4'h2][offsetY[4:0]][offsetX[4:0]] ;// wood triangle

								4'h4 : RGBout <= object_colors[4'h3][offsetY[4:0]][offsetX[4:0]] ;// wood triangle damaged

								4'h5 : RGBout <= object_colors[4'h4][offsetY[4:0]][offsetX[4:0]] ;// stone square

								4'h6 : RGBout <= object_colors[4'h5][offsetY[4:0]][offsetX[4:0]] ;// stone square damaged mid

								4'h7 : RGBout <= object_colors[4'h6][offsetY[4:0]][offsetX[4:0]] ;// stone square damaged
								
								4'h8 : RGBout <= object_colors[4'h7][offsetY[4:0]][offsetX[4:0]] ;// stone triangle

								4'h9 : RGBout <= object_colors[4'h8][offsetY[4:0]][offsetX[4:0]] ;// stone triangle damaged mid

								4'ha : RGBout <= object_colors[4'h9][offsetY[4:0]][offsetX[4:0]] ;// stone triangle damaged

								4'hb : RGBout <= object_colors[4'ha][offsetY[4:0]][offsetX[4:0]] ;// pig

								default:  RGBout <= TRANSPARENT_ENCODING ;

							endcase

						end

					end

			//--------

				HouseLoad: begin

			//--------

					if(level == 1)

					begin

						if(randomPig_LVL[8] == 1)

							MazeBitMapMask  <=  MazeLVL1B;  //  insert level 1

						else

							MazeBitMapMask  <=  MazeLVL1A;

					end

					else if(level == 2)

					begin

						if(randomPig_LVL[7] == 1)

							MazeBitMapMask  <=  MazeLVL2B;  //  insert level 2

						else

							MazeBitMapMask  <=  MazeLVL2A;

					end

					else if(level == 3)

					begin

						if(randomPig_LVL[6] == 1)

							MazeBitMapMask  <=  MazeLVL3B;  //  insert level 3

						else

							MazeBitMapMask  <=  MazeLVL3A;

					end

					levelFlag <= 1;

					SM_Motion <= PigDamageLoad;

                             

               end //HouseLoad End

                                            

			//--------

				PigDamageLoad: begin

			//--------

					if(level == 1) begin

						if(randomPig_LVL[0] == 1 && randomPig_LVL[8] == 0) //level 1 A, bottom position
						
						begin

								MazeBitMapMask[12][12] <= 4'hb;
								pigLocationX <= 12*32;
								pigLocationY <= 12*32;
						end


						else if(randomPig_LVL[0] == 0 && randomPig_LVL[8] == 0) //level 1 A, top position
						
						begin

								MazeBitMapMask[10][12] <= 4'hb;
								pigLocationX <= 12*32;
								pigLocationY <= 10*32;
								
						end


						else if(randomPig_LVL[0] == 1 && randomPig_LVL[8] == 1) //level 1 B, right position
						
						begin

								MazeBitMapMask[12][13] <= 4'hb;
								pigLocationX <= 13*32;
								pigLocationY <= 12*32;
								
						end


						else if(randomPig_LVL[0] == 0 && randomPig_LVL[8] == 1) //level 1 B, left position
						
						begin

								MazeBitMapMask[12][11] <= 4'hb;
								pigLocationX <= 11*32;
								pigLocationY <= 12*32;
								
						end


						if(randomPig_LVL[8] == 1) begin //  insert level 1B damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[10][8] <= MazeBitMapMask[10][8] + 4'h1; //block 1

								if(randomHouse[1] == 1)

										MazeBitMapMask[11][8] <= MazeBitMapMask[11][8] + 4'h1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[12][8] <= MazeBitMapMask[12][8] + 4'h1; //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 4'h1; //block 4

								if(randomHouse[4] == 1)

										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 4'h1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 4'h1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[12][10] <= MazeBitMapMask[12][10] + 4'h1; //block 7

								if(randomHouse[7] == 1)
								
										MazeBitMapMask[11][14] <= MazeBitMapMask[11][14] + 4'h1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[11][10] <= MazeBitMapMask[11][10] + 4'h1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[12][12] <= MazeBitMapMask[12][12] + 4'h1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[12][14] <= MazeBitMapMask[12][14] + 4'h1; //block 11

								end

                                                           

						else begin //insert level 1A damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[8][11] <= MazeBitMapMask[8][11] + 4'h1; //block 1

								if(randomHouse[1] == 1)

										MazeBitMapMask[8][12] <= MazeBitMapMask[8][12] + 4'h1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[8][13] <= MazeBitMapMask[8][13] + 4'h1; //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[9][11] <= MazeBitMapMask[9][11] + 4'h1; //block 4

								if(randomHouse[4] == 1)

										MazeBitMapMask[9][12] <= MazeBitMapMask[9][12] + 4'h1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[9][13] <= MazeBitMapMask[9][13] + 4'h1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[10][11] <= MazeBitMapMask[10][11] + 4'h1; //block 7

								if(randomHouse[7] == 1)

										MazeBitMapMask[10][13] <= MazeBitMapMask[10][13] + 4'h1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[11][9] <= MazeBitMapMask[11][9] + 4'h1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 4'h1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 4'h1; //block 11
										
								if(randomHouse[11] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 4'h1; //block 12

								if(randomHouse[12] == 1)

										MazeBitMapMask[12][9] <= MazeBitMapMask[12][9] + 4'h1; //block 13

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][11] <= MazeBitMapMask[12][11] + 4'h1; //block 14

								if(randomHouse[14] == 1)

										MazeBitMapMask[12][13] <= MazeBitMapMask[12][13] + 4'h1; //block 15

								end

                                                                          

					end //level1 end

                                                           

					if(level == 2) begin

                  if(randomPig_LVL[1] == 1 && randomPig_LVL[7] == 0)  //level 2 A, bottom position
						
						begin
								if(randomPig_LVL[2] == 1) //level 2, left poisition
								begin
									MazeBitMapMask[12][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 12*32;
								end
									
								else //level 2, right poisition
								begin
									MazeBitMapMask[12][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 12*32;
								end
								
						end


						else if(randomPig_LVL[1] == 0 && randomPig_LVL[7] == 0)  //level 2 A, top position
						
						begin
								if(randomPig_LVL[2] == 1) //level 2, left poisition
								begin	
									MazeBitMapMask[10][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 10*32;
								end
								
								else //level 2, right poisition
								begin	
									MazeBitMapMask[10][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 10*32;
								end
								
						end


						else if(randomPig_LVL[1] == 1 && randomPig_LVL[7] == 1)  //level 2 B, bottom position
						
						begin
								if(randomPig_LVL[2] == 1) //level 2, left poisition
								begin	
									MazeBitMapMask[12][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 12*32;
								end
									
								else //level 2, right poisition
								begin
									MazeBitMapMask[12][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 12*32;
								end
								
						end

						else if(randomPig_LVL[1] == 0 && randomPig_LVL[7] == 1)  //level 2 B, top position
						
						begin
								if(randomPig_LVL[2] == 1) //level 2, left poisition
								begin	
									MazeBitMapMask[10][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 10*32;
								end
								
								else //level 2, right poisition
								begin	
									MazeBitMapMask[10][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 10*32;
								end
								
						end
						

						if(randomPig_LVL[7] == 1) begin //  insert level 2B damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[8][11] <= MazeBitMapMask[8][11] + 1; //block 1

								if(randomHouse[1] == 1)

										MazeBitMapMask[9][7] <= MazeBitMapMask[9][7] + 1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[9][9] <= MazeBitMapMask[9][9] + 1;       //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[9][10] <= MazeBitMapMask[9][10] + 1; //block 4

								if(randomHouse[4] == 1)
										
										MazeBitMapMask[9][11] <= MazeBitMapMask[9][11] + 1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[9][12] <= MazeBitMapMask[9][12] + 1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[9][13] <= MazeBitMapMask[9][13] + 1; //block 7

								if(randomHouse[7] == 1)

										MazeBitMapMask[10][7] <= MazeBitMapMask[10][7] + 1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[10][9] <= MazeBitMapMask[10][9] + 1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[10][11] <= MazeBitMapMask[10][11] + 1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][7] <= MazeBitMapMask[11][7] + 1; //block 11

								if(randomHouse[11] == 1)

										MazeBitMapMask[11][9] <= MazeBitMapMask[11][9] + 1; //block 12

								if(randomHouse[12] == 1)

										MazeBitMapMask[11][10] <= MazeBitMapMask[11][10] + 1; //block 13

								if(randomHouse[13] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 1; //block 14

								if(randomHouse[14] == 1)

										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 1; //block 15

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 1; //block 16

								if(randomHouse[11] == 1)

										MazeBitMapMask[12][7] <= MazeBitMapMask[12][7] + 1; //block 17

								if(randomHouse[12] == 1)

										MazeBitMapMask[12][9] <= MazeBitMapMask[12][9] + 1; //block 18

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][13] <= MazeBitMapMask[12][13] + 1; //block 19

								end
								

						else begin //insert level 2A damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[8][11] <= MazeBitMapMask[8][11] + 1; //block 1

								if(randomHouse[1] == 1)
										
										MazeBitMapMask[8][12] <= MazeBitMapMask[8][12] + 1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[8][13] <= MazeBitMapMask[8][13] + 1;    //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[9][11] <= MazeBitMapMask[9][11] + 1; //block 4
										
								if(randomHouse[4] == 1)

										MazeBitMapMask[9][12] <= MazeBitMapMask[9][12] + 1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[9][13] <= MazeBitMapMask[9][13] + 1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[10][7] <= MazeBitMapMask[10][7] + 1; //block 7

								if(randomHouse[7] == 1)

										MazeBitMapMask[10][11] <= MazeBitMapMask[10][11] + 1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[10][13] <= MazeBitMapMask[10][13] + 1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[11][7] <= MazeBitMapMask[11][7] + 1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][9] <= MazeBitMapMask[11][9] + 1; //block 11
								
								if(randomHouse[11] == 1)

										MazeBitMapMask[11][10] <= MazeBitMapMask[11][10] + 1; //block 12

								if(randomHouse[12] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 1; //block 13

								if(randomHouse[13] == 1)

										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 1; //block 14
										
								if(randomHouse[14] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 1; //block 15

								if(randomHouse[10] == 1)

										MazeBitMapMask[12][7] <= MazeBitMapMask[12][7] + 1; //block 16

								if(randomHouse[11] == 1)

										MazeBitMapMask[12][9] <= MazeBitMapMask[12][9] + 1; //block 17

								if(randomHouse[12] == 1)

										MazeBitMapMask[12][11] <= MazeBitMapMask[12][11] + 1; //block 18

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][13] <= MazeBitMapMask[12][13] + 1; //block 19

								end


					end //end of level 2


					if(level == 3) begin

						if(randomPig_LVL[1] == 1 && randomPig_LVL[6] == 0)  //level 3 A, bottom position
						
						begin
								if(randomPig_LVL[2] == 1) //level 3, left poisition
								begin	
									MazeBitMapMask[12][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 12*32;
								end
								
								else //level 3, right poisition
								begin	
									MazeBitMapMask[12][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 12*32;
								end
								
						end


						else if(randomPig_LVL[1] == 0 && randomPig_LVL[6] == 0)  //level 3 A, top position
						
						begin
								if(randomPig_LVL[2] == 1) //level 3, left poisition
								begin	
									MazeBitMapMask[10][11] <= 4'hb;
									pigLocationX <= 11*32;
									pigLocationY <= 10*32;
								end
								
								else //level 3, right poisition
								begin	
									MazeBitMapMask[10][11] <= 4'hb;
									pigLocationX <= 11*32;
									pigLocationY <= 10*32;
								end
								
						end


						else if(randomPig_LVL[1] == 1 && randomPig_LVL[6] == 1)  //level 3 B, bottom position
						
						begin
								if(randomPig_LVL[2] == 1) //level 3, left poisition
								begin	
									MazeBitMapMask[12][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 12*32;
								end
								
								else //level 3, right poisition
								begin	
									MazeBitMapMask[12][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 12*32;
								end
								
						end

						else if(randomPig_LVL[1] == 0 && randomPig_LVL[6] == 1)  //level 3 B, top position
						
						begin
								if(randomPig_LVL[2] == 1) //level 3, left poisition
								begin	
									MazeBitMapMask[10][10] <= 4'hb;
									pigLocationX <= 10*32;
									pigLocationY <= 10*32;
								end
								
								else //level 3, right poisition
								begin	
									MazeBitMapMask[10][12] <= 4'hb;
									pigLocationX <= 12*32;
									pigLocationY <= 10*32;
								end
						end
						

						if(randomPig_LVL[6] == 1) begin //  insert level 3B damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[8][11] <= MazeBitMapMask[8][11] + 1; //block 1

								if(randomHouse[1] == 1)

										MazeBitMapMask[8][12] <= MazeBitMapMask[8][12] + 1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[8][13] <= MazeBitMapMask[8][13] + 1;    //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[9][9] <= MazeBitMapMask[9][9] + 1; //block 4

								if(randomHouse[4] == 1)

										MazeBitMapMask[9][11] <= MazeBitMapMask[9][11] + 1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[9][12] <= MazeBitMapMask[9][12] + 1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[9][13] <= MazeBitMapMask[9][13] + 1; //block 7

								if(randomHouse[7] == 1)

										MazeBitMapMask[10][7] <= MazeBitMapMask[10][7] + 1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[10][9] <= MazeBitMapMask[10][9] + 1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[10][11] <= MazeBitMapMask[10][11] + 1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[10][13] <= MazeBitMapMask[10][13] + 1; //block 11

								if(randomHouse[11] == 1)

										MazeBitMapMask[11][7] <= MazeBitMapMask[11][7] + 1; //block 12
										
								if(randomHouse[11] == 1)

										MazeBitMapMask[11][9] <= MazeBitMapMask[11][9] + 1; //block 13

								if(randomHouse[12] == 1)

										MazeBitMapMask[11][10] <= MazeBitMapMask[11][10] + 1; //block 14

								if(randomHouse[13] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 1; //block 15

								if(randomHouse[14] == 1)
								
										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 1; //block 16

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 1; //block 17

								if(randomHouse[11] == 1)

										MazeBitMapMask[12][7] <= MazeBitMapMask[12][7] + 1; //block 18

								if(randomHouse[12] == 1)

										MazeBitMapMask[12][9] <= MazeBitMapMask[12][9] + 1; //block 19

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][11] <= MazeBitMapMask[12][11] + 1; //block 20

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][13] <= MazeBitMapMask[12][13] + 1; //block 21

								end

                                                                          

                                                           

						else begin //insert level 3A damage

								if(randomHouse[0] == 1)

										MazeBitMapMask[8][10] <= MazeBitMapMask[8][10] + 1; //block 1

								if(randomHouse[1] == 1)

										MazeBitMapMask[8][11] <= MazeBitMapMask[8][11] + 1; //block 2

								if(randomHouse[2] == 1)

										MazeBitMapMask[8][12] <= MazeBitMapMask[8][12] + 1;    //block 3

								if(randomHouse[3] == 1)

										MazeBitMapMask[9][10] <= MazeBitMapMask[9][10] + 1; //block 4

								if(randomHouse[4] == 1)

										MazeBitMapMask[9][11] <= MazeBitMapMask[9][11] + 1; //block 5

								if(randomHouse[5] == 1)

										MazeBitMapMask[9][12] <= MazeBitMapMask[9][12] + 1; //block 6

								if(randomHouse[6] == 1)

										MazeBitMapMask[10][7] <= MazeBitMapMask[10][7] + 1; //block 7
								
								if(randomHouse[7] == 1)

										MazeBitMapMask[10][9] <= MazeBitMapMask[10][9] + 1; //block 8

								if(randomHouse[8] == 1)

										MazeBitMapMask[10][10] <= MazeBitMapMask[10][10] + 1; //block 9

								if(randomHouse[9] == 1)

										MazeBitMapMask[10][12] <= MazeBitMapMask[10][12] + 1; //block 10

								if(randomHouse[10] == 1)

										MazeBitMapMask[10][13] <= MazeBitMapMask[10][13] + 1; //block 11

								if(randomHouse[11] == 1)

										MazeBitMapMask[11][7] <= MazeBitMapMask[11][7] + 1; //block 12

								if(randomHouse[11] == 1)
								
										MazeBitMapMask[11][9] <= MazeBitMapMask[11][9] + 1; //block 13
										
								if(randomHouse[12] == 1)

										MazeBitMapMask[11][10] <= MazeBitMapMask[11][10] + 1; //block 14

								if(randomHouse[13] == 1)

										MazeBitMapMask[11][11] <= MazeBitMapMask[11][11] + 1; //block 15

								if(randomHouse[14] == 1)

										MazeBitMapMask[11][12] <= MazeBitMapMask[11][12] + 1; //block 16

								if(randomHouse[10] == 1)

										MazeBitMapMask[11][13] <= MazeBitMapMask[11][13] + 1; //block 17

								if(randomHouse[11] == 1)

										MazeBitMapMask[12][7] <= MazeBitMapMask[12][7] + 1; //block 18
								if(randomHouse[12] == 1)

										MazeBitMapMask[12][9] <= MazeBitMapMask[12][9] + 1; //block 19

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][11] <= MazeBitMapMask[12][11] + 1; //block 20

								if(randomHouse[13] == 1)

										MazeBitMapMask[12][13] <= MazeBitMapMask[12][13] + 1; //block 21

								end

                                            

					end //end of level 3

                                            

					SM_Motion <= Idle;

                                                           

				end//PigDamageLoad End
				
				
				//--------

				WinningScreen: begin //WinningScreen Start

				//--------
						enterKey_D <= enterKey;
						if(enterKey && !enterKey_D) begin
							SM_Motion <= Idle;
							level1Vic <= 0;
							level2Vic <= 0;
							level3Vic <= 0;
							levelFlag <= 0;
						end
				
				end //WinningScreen End

      endcase

	end 
end
 

//==----------------------------------------------------------------------------------------------------------------=

// decide if to draw the pixel or not

assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap

assign fire = ( (MazeBitMapMask[randomX][randomY] == 4'h1) ||   

                (MazeBitMapMask[randomX][randomY] == 4'h2) ||

                (MazeBitMapMask[randomX][randomY] == 4'h3) ||

                (MazeBitMapMask[randomX][randomY] == 4'h4) ||

                (MazeBitMapMask[randomX][randomY] == 4'h5)  ) ? 1'b1 : 1'b0;

 

  

endmodule